// reloj.v

// Generated using ACDS version 22.1 915

`timescale 1 ps / 1 ps
module reloj (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

endmodule
